module overlap_243bit(p0,p1,p2,p3,p4,p5,y);
input [160:0] p0,p1,p2,p3,p4,p5;
output [484:0] y;

assign y[80:0] = p0[80:0];
assign y[160:81] = p0[160:81]^p0[79:0]^p1[79:0]^p2[79:0];
assign y[161] = p0[80]^p1[80]^p2[80];
assign y[241:162] = p0[160:81]^p1[160:81]^p2[160:81]^p0[79:0]^p1[79:0]^p3[79:0]^p4[79:0];
assign y[242] = p0[80]^p1[80]^p3[80]^p4[80];
assign y[322:243] = p0[160:81]^p1[160:81]^p3[160:81]^p4[160:81]^p1[79:0]^p3[79:0]^p5[79:0];
assign y[323] = p1[80]^p5[80]^p3[80];
assign y[403:324] = p1[160:81]^p5[160:81]^p3[160:81]^p3[79:0];
assign y[484:404] = p3[160:80];

endmodule
