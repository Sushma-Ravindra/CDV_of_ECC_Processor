module overlap_81bit(p0,p1,p2,p3,p4,p5,y);
input [52:0] p0,p1,p2,p3,p4,p5;
output [160:0] y;

assign y[26:0] = p0[26:0];
assign y[52:27] = p0[52:27]^p0[25:0]^p1[25:0]^p2[25:0];
assign y[53] = p0[26]^p1[26]^p2[26];
assign y[79:54] = p0[52:27]^p1[52:27]^p2[52:27]^p0[25:0]^p1[25:0]^p3[25:0]^p4[25:0];
assign y[80] = p0[26]^p1[26]^p3[26]^p4[26];
assign y[106:81] = p0[52:27]^p1[52:27]^p3[52:27]^p4[52:27]^p1[25:0]^p3[25:0]^p5[25:0];
assign y[107] = p1[26]^p5[26]^p3[26];
assign y[133:108] = p1[52:27]^p5[52:27]^p3[52:27]^p3[25:0];
assign y[160:134] = p3[52:26];

endmodule
